library verilog;
use verilog.vl_types.all;
entity uart_test_pkg is
end uart_test_pkg;
